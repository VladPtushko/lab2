library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use ieee.std_logic_unsigned.all;

entity sin_lut is
    port (
        address_a		: IN STD_LOGIC_VECTOR (7 DOWNTO 0) := (others => '0') ;
		address_b		: IN STD_LOGIC_VECTOR (7 DOWNTO 0) := (others => '0') ;
		clock		: IN STD_LOGIC  := '1';
		q_a		: OUT STD_LOGIC_VECTOR (8 DOWNTO 0) := (others => '0');
		q_b		: OUT STD_LOGIC_VECTOR (8 DOWNTO 0) := (others => '0')
    );
end entity sin_lut;

architecture a_sin_lut of sin_lut is
    TYPE int_array is ARRAY (natural range <>) of integer;            -- int_array type declaration

    CONSTANT lut : int_array := (                                     -- Look up table cells/arrays
        0,
        3,
        6,
        9,
        13,
        16,
        19,
        22,
        25,
        28,
        31,
        34,
        38,
        41,
        44,
        47,
        50,
        53,
        56,
        59,
        63,
        66,
        69,
        72,
        75,
        78,
        81,
        84,
        87,
        90,
        94,
        97,
        100,
        103,
        106,
        109,
        112,
        115,
        118,
        121,
        124,
        127,
        130,
        133,
        136,
        139,
        142,
        145,
        148,
        151,
        154,
        157,
        160,
        163,
        166,
        169,
        172,
        175,
        178,
        181,
        184,
        187,
        190,
        193,
        196,
        198,
        201,
        204,
        207,
        210,
        213,
        216,
        218,
        221,
        224,
        227,
        230,
        233,
        235,
        238,
        241,
        244,
        246,
        249,
        252,
        255,
        257,
        260,
        263,
        265,
        268,
        271,
        273,
        276,
        279,
        281,
        284,
        286,
        289,
        292,
        294,
        297,
        299,
        302,
        304,
        307,
        309,
        312,
        314,
        317,
        319,
        322,
        324,
        327,
        329,
        331,
        334,
        336,
        338,
        341,
        343,
        345,
        348,
        350,
        352,
        355,
        357,
        359,
        361,
        364,
        366,
        368,
        370,
        372,
        374,
        377,
        379,
        381,
        383,
        385,
        387,
        389,
        391,
        393,
        395,
        397,
        399,
        401,
        403,
        405,
        407,
        409,
        410,
        412,
        414,
        416,
        418,
        420,
        421,
        423,
        425,
        427,
        428,
        430,
        432,
        433,
        435,
        437,
        438,
        440,
        441,
        443,
        445,
        446,
        448,
        449,
        451,
        452,
        454,
        455,
        456,
        458,
        459,
        461,
        462,
        463,
        465,
        466,
        467,
        468,
        470,
        471,
        472,
        473,
        474,
        476,
        477,
        478,
        479,
        480,
        481,
        482,
        483,
        484,
        485,
        486,
        487,
        488,
        489,
        490,
        491,
        492,
        492,
        493,
        494,
        495,
        496,
        496,
        497,
        498,
        499,
        499,
        500,
        501,
        501,
        502,
        502,
        503,
        503,
        504,
        505,
        505,
        505,
        506,
        506,
        507,
        507,
        508,
        508,
        508,
        509,
        509,
        509,
        509,
        510,
        510,
        510,
        510,
        510,
        511,
        511,
        511,
        511,
        511,
        511,
        511
    );

    SIGNAL lut_address_index_a : integer range 0 to 255;
    SIGNAL lut_address_index_b : integer range 0 to 255;

begin
    lut_address_index_a <= CONV_INTEGER(unsigned(address_a));           
    q_a <= std_logic_vector(CONV_UNSIGNED(lut(lut_address_index_a), q_a'length));  
    
    lut_address_index_b <= CONV_INTEGER(unsigned(address_b));           
    q_b <= std_logic_vector(CONV_UNSIGNED(lut(lut_address_index_b), q_b'length)); 
end architecture;